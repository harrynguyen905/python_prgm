module test ()


input
output

endmodule

