module test ()
endmodule

